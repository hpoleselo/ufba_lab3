library verilog;
use verilog.vl_types.all;
entity interfaceCC_vlg_vec_tst is
end interfaceCC_vlg_vec_tst;
